module Segment7(num, segs);
input [3:0] num ; //the hex digit to be displayed
output [6:0] segs ; //actual LED segments
reg [6:0] segs ;
always @ (num)
begin
case (num)
4'h0: segs = 7'b1000000;
4'h1: segs = 7'b1111001;
4'h2: segs = 7'b0100100;
4'h3: segs = 7'b0110000;
4'h4: segs = 7'b0011001;
4'h5: segs = 7'b0010010;
4'h6: segs = 7'b0000010;
4'h7: segs = 7'b1111000;
4'h8: segs = 7'b0000000;
4'h9: segs = 7'b0010000;
4'ha: segs = 7'b0001000;
4'hb: segs = 7'b0000011;
4'hc: segs = 7'b1000110;
4'hd: segs = 7'b0100001;
4'he: segs = 7'b0000110;
4'hf: segs = 7'b0001110;
default segs = 7'b1111111;
endcase
end
endmodule